module pgMatricula();

  logic        clk;
  logic        reset;

  logic [31:0] WriteData, DataAdr;
  logic        MemWrite;

  // instantiate device to be tested
  top dut(clk, reset, WriteData, DataAdr, MemWrite);
  
  // initialize test
  initial
    begin
      reset <= 1; # 22; reset <= 0;
	//reset <= 0;
    end

  // generate clock to sequence tests
  always
    begin
      clk <= 1; # 5; clk <= 0; # 5;
    end

  // check results
  always @(negedge clk)
    begin
      if(MemWrite) begin
        if(WriteData === 166912) begin
          $display("Simulation succeeded");
          $stop;
        //end else if (WriteData !== 1 & WriteData !== 2 & WriteData !== 3 & WriteData !== 5) begin //| WriteData !== 3 | WriteData !== 5 | WriteData !== 5
        //  $display("Simulation failed");
        //  $stop;
        end
      end
    end
endmodule